-------------------------------------------------------------------------------
-- Title      : DLX_top
-- Project    : 
-------------------------------------------------------------------------------
-- File       : DLX_top.vhd
-- Author     :   <michel agoyan@ROU13572>
-- Company    : 
-- Created    : 2015-11-25
-- Last update: 2019-08-23
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: DLX data path + control path
-------------------------------------------------------------------------------
-- Copyright (c) 2019 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2015-11-25  1.0      michel agoyan   Created
-- 2019-08-21  1.1      Olivier potin   Modified to implement RISCV Monocycle
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
library rtl_core;
use rtl_core.RV32I_components.all;
use rtl_core.RV32I_constants.all;

library rtl_tracer;

entity RV32I_Monocycle_top is

  generic (
    rom_init_filename: string:="rom.hex";
	ram_init_filename: string:=""; 
	TLEN : POSITIVE);

  port (
    clk_i        : in std_logic;
	resetn_i     : in std_logic;
	enable_tracer_i : in std_logic;
	trace_o		 : out std_logic_vector((TLEN*8)-1 downto 0);
	trace_length_o : out NATURAL range 0 to (TLEN-1);
	trace_emitted_o : out std_logic;
	PeriphAddr_o : out std_logic_vector(31 downto 0); -- Periph address
    PeriphData_o : out std_logic_vector(31 downto 0); -- Periph word
    PeriphWe_o   : out std_logic); -- set when Periph word is valid

end entity RV32I_Monocycle_top;

architecture RV32I_Monocycle_top_architecture of RV32I_Monocycle_top is
-- component declaration
component RV32I_TraceEncoder is
    generic (TLEN : POSITIVE);
    port (  clock_i : in std_logic;
            resetb_i : in std_logic;
            enable_i : in std_logic;
            exception_i : in std_logic; -- an exception occurs
            iaddr_i : in std_logic_vector(IADDRESS_WIDTH_P-1 downto 0);   -- next instruction address
            instr_i : in std_logic_vector(INSTR_WIDTH_P-1 downto 0);        -- current instruction
            ecause_i : in std_logic_vector(MCAUSE_WIDTH_P-1 downto 0);
            tval_i : in std_logic_vector(IADDRESS_WIDTH_P-1 downto 0);
            priv_i : in std_logic_vector(PRIVILEGE_WIDTH_P-1 downto 0);   -- fixed as user privilege for us
            trace_o : out std_logic_vector((TLEN*8)-1 downto 0);
            trace_length_o : out NATURAL range 0 to (TLEN-1);
	        trace_emitted_o : out std_logic);
end component;

-- RV32 current instruction (i.e from datapath to control path) 
-- see Patterson & Hennessy page  257 for global sheme
signal Instruction_s : std_logic_vector(31 downto 0);
-- outputs signal generated by controler (i.e from controlpath to datapath)
-- see patterson and Hennessy page 256
signal IAddress_s : std_logic_vector(31 downto 0);  -- current instruction address 
signal MemRead_s : std_logic;
signal MemWrite_s : std_logic;
signal MemSelectData_s : std_logic_vector(2 downto 0);
signal RegWrite_s : std_logic; 
signal ALUSrc1_s : std_logic_vector(1 downto 0);
signal ALUSrc2_s : std_logic_vector(0 downto 0);
signal ALU_zero_s : std_logic;
signal ALU_lt_s : std_logic;
signal ALU_ltu_s : std_logic;
signal ALUControl_s : std_logic_vector(3 downto 0);
signal WB_select_s : std_logic_vector(1 downto 0);
signal PC_select_s : std_logic_vector(1 downto 0);
signal exception_s : std_logic;
signal unknown_instr_s : std_logic;
signal tval_s : std_logic_vector(IADDRESS_WIDTH_P-1 downto 0);
signal mcause_s : std_logic_vector(MCAUSE_WIDTH_P-1 downto 0);
begin  -- architecture RV32I_Monocycle_top_architecture

  RV32I_Monocycle_controlpath_1 : RV32I_Monocycle_controlpath
    port map (
	Instruction_i	=> Instruction_s,
	ALU_zero_i	=> ALU_zero_s,
	ALU_lt_i	=> ALU_lt_s,	
	ALU_ltu_i	=> ALU_ltu_s,	
	exception_i => exception_s,
	unknown_instr_o => unknown_instr_s,	
	PC_select_o	=> PC_select_s,	
	ALUSrc1_o	=> ALUSrc1_s,
	ALUSrc2_o	=> ALUSrc2_s,
	ALUControl_o	=> ALUControl_s,
	MemWrite_o	=> MemWrite_s,
	MemRead_o	=> MemRead_s,
	MemSelectData_o => MemSelectData_s,
	WB_select_o	=> WB_select_s,
	RegWrite_o	=> RegWrite_s);

  RV32I_Monocycle_datapath_1 : RV32I_Monocycle_datapath
    generic map (
	rom_init_filename => rom_init_filename,
	ram_init_filename => ram_init_filename
    ) port map (
	clk_i		=> clk_i,
	resetn_i	=> resetn_i,
	IAddress_o	=> IAddress_s,
	Instruction_o	=> Instruction_s,
	ALU_zero_o	=> ALU_zero_s,
	ALU_lt_o	=> ALU_lt_s,	
	ALU_ltu_o	=> ALU_ltu_s,	
	PC_select_i	=> PC_select_s,	
	ALUSrc1_i	=> ALUSrc1_s,
	ALUSrc2_i	=> ALUSrc2_s,
	ALUControl_i	=> ALUControl_s,
	MemWrite_i	=> MemWrite_s,
	MemRead_i	=> MemRead_s,
	MemSelectData_i => MemSelectData_s,
	WB_select_i	=> WB_select_s,
	RegWrite_i	=> RegWrite_s,
	unknown_instr_i => unknown_instr_s,	
	exception_o 	=> exception_s,
	tval_o 		=> tval_s,
	mcause_o 	=> mcause_s,
	PeriphAddr_o	=> PeriphAddr_o,
	PeriphData_o	=> PeriphData_o,
	PeriphWe_o	=> PeriphWe_o);

	UTracer: RV32I_TraceEncoder 
	generic map (TLEN => TLEN)		
	port map (  
		clock_i => clk_i,
		resetb_i => resetn_i,
		enable_i => enable_tracer_i,
		exception_i => exception_s,
		iaddr_i => IAddress_s, 
		instr_i => Instruction_s,
		ecause_i => mcause_s,
		tval_i => tval_s,
		priv_i => "00",
		trace_o => trace_o,
		trace_length_o => trace_length_o,
		trace_emitted_o => trace_emitted_o);
	
end architecture RV32I_Monocycle_top_architecture;

-------------------------------------------------------------------------------
-- Title      : DLX_top
-- Project    : 
-------------------------------------------------------------------------------
-- File       : DLX_top.vhd
-- Author     :   <michel agoyan@ROU13572>
-- Company    : 
-- Created    : 2015-11-25
-- Last update: 2019-08-23
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: DLX data path + control path
-------------------------------------------------------------------------------
-- Copyright (c) 2019 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2015-11-25  1.0      michel agoyan   Created
-- 2019-08-21  1.1      Olivier potin   Modified to implement RISCV Pipelined
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use work.RV32I_components.all;

entity RV32I_Pipelined_top is

  port (
    clk_i    : in std_logic;
    resetn_i : in std_logic);

end entity RV32I_Pipelined_top;

architecture RV32I_Pipelined_top_architecture of RV32I_Pipelined_top is
-- RV32 instructions in stages (i.e from datapath to control path) 
-- see Patterson & Hennessy page 294 for global sheme
signal Instruction_IFID_s : std_logic_vector(31 downto 0);
signal Instruction_IDEX_s : std_logic_vector(25 downto 0);
signal Instruction_EXMEM_s : std_logic_vector(14 downto 0);
signal Instruction_MEMWB_s : std_logic_vector(4 downto 0);
-- outputs signal generated by controler (i.e from controlpath to datapath)
-- see patterson and Hennessy page 294
signal MemRead_s : std_logic;
signal MemWrite_s : std_logic;
signal RegWrite_s : std_logic; 
signal ALUSrc1_s : std_logic_vector(1 downto 0);
signal ALUSrc2_s : std_logic_vector(0 downto 0);
signal ALU_zero_s : std_logic;
signal ALU_lt_s : std_logic;
signal ALUControl_s : std_logic_vector(3 downto 0);
Signal ForwardA_s : std_logic_vector(1 downto 0);
Signal ForwardB_s : std_logic_vector(1 downto 0);
signal WB_select_s : std_logic_vector(1 downto 0);
signal PC_select_s : std_logic_vector(1 downto 0);
signal PCWrite_s : std_logic;
signal IFIDWrite_s : std_logic;
begin  -- architecture RV32I_Pipelined_top_architecture

  RV32I_Pipelined_controlpath_1 : RV32I_Pipelined_controlpath
    port map (
	clk_i 		=> clk_i,
	resetn_i 	=> resetn_i,
	Instruction_IFID_i	=> Instruction_IFID_s,
	Instruction_IDEX_i	=> Instruction_IDEX_s,
	Instruction_EXMEM_i	=> Instruction_EXMEM_s,
	Instruction_MEMWB_i	=> Instruction_MEMWB_s,
	ALU_zero_i	=> ALU_zero_s,
	ALU_lt_i	=> ALU_lt_s,	
	PC_select_o	=> PC_select_s,	
	ALUSrc1_o	=> ALUSrc1_s,
	ALUSrc2_o	=> ALUSrc2_s,
	ALUControl_o	=> ALUControl_s,
	ForwardA_o	=> ForwardA_s,
	ForwardB_o	=> ForwardB_s,
	MemWrite_o	=> MemWrite_s,
	MemRead_o	=> MemRead_s,
	WB_select_o	=> WB_select_s,
	RegWrite_o	=> RegWrite_s,
	PCWrite_o	=> PCWrite_s,
	IFIDWrite_o	=> IFIDWrite_s);	

  RV32I_Pipelined_datapath_1 : RV32I_Pipelined_datapath
    port map (
	clk_i		=> clk_i,
	resetn_i	=> resetn_i,
	Instruction_IFID_o	=> Instruction_IFID_s,
	Instruction_IDEX_o	=> Instruction_IDEX_s,
	Instruction_EXMEM_o	=> Instruction_EXMEM_s,
	Instruction_MEMWB_o	=> Instruction_MEMWB_s,
	ALU_zero_o	=> ALU_zero_s,
	ALU_lt_o	=> ALU_lt_s,	
	PC_select_i	=> PC_select_s,	
	ALUSrc1_i	=> ALUSrc1_s,
	ALUSrc2_i	=> ALUSrc2_s,
	ALUControl_i	=> ALUControl_s,
	ForwardA_i	=> ForwardA_s,
	ForwardB_i	=> ForwardB_s,
	MemWrite_i	=> MemWrite_s,
	MemRead_i	=> MemRead_s,
	WB_select_i	=> WB_select_s,
	RegWrite_i	=> RegWrite_s,	
	PCWrite_i	=> PCWrite_s,
	IFIDWrite_i	=> IFIDWrite_s);

end architecture RV32I_Pipelined_top_architecture;
